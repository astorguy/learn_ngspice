* Voltage Divider Circuit Example
V1 in 0 DC 10V
R1 in out 1k
R2 out 0 2k

* Analysis Command: Calculate DC Operating Point
.op
.end
